library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- La pista rotada para evitar utilizar una memoria y gestionar los accesos
package not_Mapatrack_pkg is

  type memoracetrack is array (natural range<>) of
       std_logic_vector(32-1 downto 0);
  constant not_pista : memoracetrack := (
       "00000000000000000000000000000000",
       "00000000000000000000000000000000",
       "00000000000000000000000000000000",
       "00000000000000000000000000000000",
       "00000000000000000000000000000000",
       "00011111111111111111111111111000",
       "00011111111111111111111111111000",
       "00001111111111111111000011111000",
       "00000011111111111111100111111000",
       "00000011111111111111111111111000",
       "00000001111111111111111111111000",
       "00000011111111111111111111111000",
       "00001111111111111111111111111000",
       "00011111111111111111111111111000",
       "00011111100111111111111111111111",
       "00011111100111111111111111111111",
       "00011111100111111111111111111111",
       "00011111111111111111111111111111",
       "00011111111111111101111111111111",
       "00011111111111111000111111111000",
       "00011111111111111100111111111000",
       "00011111111111111111111111111000",
       "00011111111111111111111111110000",
       "00011111111111111111111111100000",
       "00011111111111111111111110000000",
       "00011111100111111111111111100000",
       "00011111100011111111111111110000",
       "00011111110011111111111111111000",
       "00011111111111111111111111111000",
       "00000000000000000001111100000000"
        );

end not_Mapatrack_pkg;

